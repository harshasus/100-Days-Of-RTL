`timescale 1ns / 1ps
module inv(input a,output b);
assign b=~a;
endmodule
